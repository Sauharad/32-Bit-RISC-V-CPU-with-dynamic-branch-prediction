`timescale 1ns / 1ps


module UART_peripheral();



endmodule
